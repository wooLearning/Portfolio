module Window3x3_RGB888#(
	parameter DATA_W = 24,
	parameter ADDR_W = 17,
	parameter WIDTH = 480,
	parameter HEIGHT = 272,
	parameter DEPTH  = 130560
)(
	input iClk,
	input iRst,
	input iEn,

	/*for bram*/
	output oCs,
	output [ADDR_W-1 : 0] oAddr,
	input  [DATA_W-1 : 0] iPixel,

	/*next block 3x3 pixel */
	output [DATA_W-1:0] oOut0,
	output [DATA_W-1:0] oOut1,
	output [DATA_W-1:0] oOut2,
	output [DATA_W-1:0] oOut3,
	output [DATA_W-1:0] oOut4,
	output [DATA_W-1:0] oOut5,
	output [DATA_W-1:0] oOut6,
	output [DATA_W-1:0] oOut7,
	output [DATA_W-1:0] oOut8,
	output oValid
	
);

localparam IDLE = 4'd0;
localparam FIRST_ROW_FILL = 4'd1;
localparam FIRST_ROW = 4'd2;
localparam MIDDLE_ROW = 4'd3;
localparam LAST_ROW = 4'd4;
//fsm
reg [3:0] cur_state;
reg [3:0] nxt_state;
//part1
always @(posedge iClk or negedge iRst) begin
	if(!iRst) begin
		cur_state <= IDLE;
	end
	else if(iEn == 1'b1)begin
		cur_state <= nxt_state;
	end
	else begin
		cur_state <= cur_state;
	end
end

//part2
always @(*) begin
	case (cur_state)
		IDLE: begin
			if(iEn == 1'b1) nxt_state = FIRST_ROW_FILL; else nxt_state = IDLE;
		end 
		FIRST_ROW_FILL : begin
			if(rAddr_d2 == WIDTH - 1) nxt_state = FIRST_ROW; else nxt_state = FIRST_ROW_FILL;
		end
		FIRST_ROW: begin
			if(wColEnd) nxt_state = MIDDLE_ROW; else nxt_state = FIRST_ROW;
		end
		MIDDLE_ROW : begin
			if(rRowCnt == HEIGHT -2) nxt_state =LAST_ROW; else nxt_state = MIDDLE_ROW;
		end
		LAST_ROW: begin
			if(wRowEnd) nxt_state = IDLE; else nxt_state = LAST_ROW;
		end
		default:nxt_state = IDLE; 
	endcase
end

integer i;

reg [ADDR_W-1:0] rAddr;
always @(posedge iClk or negedge iRst) begin
	if(!iRst) begin
		rAddr <= 0;
	end
	else if(iEn == 1'b1)begin
		if(rAddr == (WIDTH*HEIGHT - 1)) begin
			rAddr <= 0;
		end
		else if(cur_state == IDLE) begin
			rAddr <= 0;
		end
		else begin
			rAddr <= rAddr + 1'b1;
		end
	end
	else begin
		rAddr <= rAddr;
	end
end

// 파이프라인 레지스터 (Delay용)
reg [ADDR_W -1 : 0] rAddr_d1;
reg [ADDR_W -1 : 0] rAddr_d2;
always @(posedge iClk or negedge iRst) begin
	if(!iRst) begin
		rAddr_d1 <= 0;
		rAddr_d2 <= 0;
	end
	else if(cur_state == IDLE) begin
		rAddr_d1 <= 0;
		rAddr_d2 <= 0;
	end
	else if(iEn == 1'b1) begin
		rAddr_d1 <= rAddr;
		rAddr_d2 <= rAddr_d1;
	end
end

wire wColEnd = (rColCnt == WIDTH-1);
wire wRowEnd = (rRowCnt == HEIGHT-1);

reg [$clog2(WIDTH) -1 : 0] rColCnt;

always @(posedge iClk or negedge iRst) begin
	if(!iRst) begin
		rColCnt <= 0;
	end 
	else if (wOValid && iEn == 1'b1) begin
		if (wColEnd) begin
			rColCnt <= 0;
		end
		else begin
			rColCnt <= rColCnt + 1'b1;
		end
	end
end

reg [$clog2(HEIGHT) -1 : 0] rRowCnt;
always @(posedge iClk or negedge iRst) begin
	if(!iRst) begin
		rRowCnt <= 0;
	end 
	else if (wOValid && iEn == 1'b1) begin
		if (rRowCnt == HEIGHT) begin
			rRowCnt <= 0;
		end
		else if(wColEnd) begin //timing 봐야함
			rRowCnt <= rRowCnt + 1'b1;
		end
	end
end

reg [DATA_W-1:0] rLineBuf0 [0:WIDTH-1]; 
reg [DATA_W-1:0] rLineBuf1 [0:WIDTH-1];
reg [DATA_W-1:0] rPix[0:2];
reg [1:0] rPixCnt;

always @(posedge iClk or negedge iRst) begin
	if(!iRst)begin
		for (i=0; i<WIDTH;i=i+1 ) begin
			rLineBuf0[i] <= 0;
			rLineBuf1[i] <= 0;
		end
		for(i=0;i<3;i=i+1) begin
			rPix[i] <= 0;
		end
		rPixCnt <= 0;
	end
	else if(iEn == 1'b1) begin
		case (cur_state)
			IDLE : begin
				rPixCnt <= 0;
			end
			FIRST_ROW_FILL: begin
				rLineBuf1[WIDTH-1] <= iPixel;
				for(i=WIDTH-2; i>=0; i=i-1) begin
					rLineBuf1[i] <= rLineBuf1[i+1];
				end
				rLineBuf0[WIDTH-1] <= iPixel;
				for(i=WIDTH-2; i>=0; i=i-1) begin
					rLineBuf0[i] <= rLineBuf0[i+1];
				end
			end 
			default: begin
				rPix[2] <= iPixel;
				rPix[1] <= rPix[2];
				rPix[0] <= rPix[1];
				rLineBuf1[rColCnt] <= rPix[0];
			end
		endcase
	end
end

wire wOValid = (cur_state != FIRST_ROW_FILL)&&(cur_state != IDLE)  ? 1 : 0;
reg [DATA_W-1:0] wOut[0:8];

//part3
assign wOut[0] = (cur_state == FIRST_ROW) ? 0 : 
				 (rColCnt == 0) ? 0 : rLineBuf0[rColCnt-1];
assign wOut[1] = (cur_state == FIRST_ROW) ? 0 : rLineBuf0[rColCnt];
assign wOut[2] = (cur_state == FIRST_ROW) ? 0 : rLineBuf0[rColCnt+1];

assign wOut[3] = (rColCnt == 0) ? 0 : rLineBuf1[rColCnt-1];
assign wOut[4] = rLineBuf1[rColCnt];
assign wOut[5] = rLineBuf1[rColCnt+1];

assign wOut[6] = (cur_state == LAST_ROW) ? 0 : 
				 (rColCnt == 0) ? 0 : rPix[0];
assign wOut[7] = (cur_state == LAST_ROW) ? 0 rPix[1];
assign wOut[8] = (cur_state == LAST_ROW) ? 0rPix[2];

assign oOut0 = wOut[0];
assign oOut1 = wOut[1];
assign oOut2 = wOut[2];
assign oOut3 = wOut[3];
assign oOut4 = wOut[4];
assign oOut5 = wOut[5];
assign oOut6 = wOut[6];
assign oOut7 = wOut[7];
assign oOut8 = wOut[8];
assign oValid = wOValid;

assign oCs = iEn && !((cur_state == IDLE));
assign oAddr = rAddr;
endmodule
